`timescale 1ns / 1ps
module CPU();
    
endmodule
